----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:42:34 02/25/2020 
-- Design Name: 
-- Module Name:    RF_WA_mux - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity RF_WA_mux is
    Port ( IR_15_11 : in  STD_LOGIC_VECTOR (4 downto 0);
           IR_20_16 : in  STD_LOGIC_VECTOR (4 downto 0);
			  RF_WA_MUX : in STD_LOGIC_VECTOR (1 downto 0);
           WA : out  STD_LOGIC_VECTOR (4 downto 0));
end RF_WA_mux;

architecture Behavioral of RF_WA_mux is

begin
   with RF_WA_MUX select
      WA <=    IR_15_11          when "00",
               IR_20_16          when "01",
					"11110"           when "10",
       	   	"11111"           when others;

			

end Behavioral;

